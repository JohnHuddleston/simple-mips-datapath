//////////////////////////////////////////////////////////////////////////////////
//										
// 32-bit Mux							
// 										
//////////////////////////////////////////////////////////////////////////////////

module FullMux(
	input [31:0] a, b,
	input select;
	output reg out
	);

	assign out = (select == 0?) a : b;

endmodule